library IEEE;
use IEEE.numeric_std.all;
use IEEE.std_logic_1164.all;

package TemplatePackage is
end package;

package body TemplatePackage is
end package body;
